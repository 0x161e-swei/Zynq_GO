parameter [0:7]char_rom[0:1535]={
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,// space 8'h20
8'h00,
8'h00,
8'h18,
8'h3C,
8'h3C,
8'h3C,
8'h18,
8'h18,
8'h18,
8'h00,
8'h18,
8'h18,
8'h00,
8'h00,
8'h00,
8'h00,// !
8'h00,
8'h63,
8'h63,
8'h63,
8'h22,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,// "
8'h00,
8'h00,
8'h00,
8'h36,
8'h36,
8'h7F,
8'h36,
8'h36,
8'h36,
8'h7F,
8'h36,
8'h36,
8'h00,
8'h00,
8'h00,
8'h00,// #
8'h0C,
8'h0C,
8'h3E,
8'h63,
8'h61,
8'h60,
8'h3E,
8'h03,
8'h03,
8'h43,
8'h63,
8'h3E,
8'h0C,
8'h0C,
8'h00,
8'h00,// $
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h61,
8'h63,
8'h06,
8'h0C,
8'h18,
8'h33,
8'h63,
8'h00,
8'h00,
8'h00,
8'h00,// %
8'h00,
8'h00,
8'h00,
8'h1C,
8'h36,
8'h36,
8'h1C,
8'h3B,
8'h6E,
8'h66,
8'h66,
8'h3B,
8'h00,
8'h00,
8'h00,
8'h00,// &
8'h00,
8'h30,
8'h30,
8'h30,
8'h60,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,// '
8'h00,
8'h00,
8'h0C,
8'h18,
8'h18,
8'h30,
8'h30,
8'h30,
8'h30,
8'h18,
8'h18,
8'h0C,
8'h00,
8'h00,
8'h00,
8'h00,// (
8'h00,
8'h00,
8'h18,
8'h0C,
8'h0C,
8'h06,
8'h06,
8'h06,
8'h06,
8'h0C,
8'h0C,
8'h18,
8'h00,
8'h00,
8'h00,
8'h00,// )
8'h00,
8'h00,
8'h00,
8'h00,
8'h42,
8'h66,
8'h3C,
8'hFF,
8'h3C,
8'h66,
8'h42,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,// *
8'h00,
8'h00,
8'h00,
8'h00,
8'h18,
8'h18,
8'h18,
8'hFF,
8'h18,
8'h18,
8'h18,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,// +
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h18,
8'h18,
8'h18,
8'h30,
8'h00,
8'h00,// ,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'hFF,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,// -
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h18,
8'h18,
8'h00,
8'h00,
8'h00,
8'h00,// .
8'h00,
8'h00,
8'h01,
8'h03,
8'h07,
8'h0E,
8'h1C,
8'h38,
8'h70,
8'hE0,
8'hC0,
8'h80,
8'h00,
8'h00,
8'h00,
8'h00,// / (forward slash)
8'h00,
8'h00,
8'h3E,
8'h63,
8'h63,
8'h63,
8'h6B,
8'h6B,
8'h63,
8'h63,
8'h63,
8'h3E,
8'h00,
8'h00,
8'h00,
8'h00,// 0 8'h30
8'h00,
8'h00,
8'h0C,
8'h1C,
8'h3C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h3F,
8'h00,
8'h00,
8'h00,
8'h00,// 1
8'h00,
8'h00,
8'h3E,
8'h63,
8'h03,
8'h06,
8'h0C,
8'h18,
8'h30,
8'h61,
8'h63,
8'h7F,
8'h00,
8'h00,
8'h00,
8'h00,// 2
8'h00,
8'h00,
8'h3E,
8'h63,
8'h03,
8'h03,
8'h1E,
8'h03,
8'h03,
8'h03,
8'h63,
8'h3E,
8'h00,
8'h00,
8'h00,
8'h00,// 3
8'h00,
8'h00,
8'h06,
8'h0E,
8'h1E,
8'h36,
8'h66,
8'h66,
8'h7F,
8'h06,
8'h06,
8'h0F,
8'h00,
8'h00,
8'h00,
8'h00,// 4
8'h00,
8'h00,
8'h7F,
8'h60,
8'h60,
8'h60,
8'h7E,
8'h03,
8'h03,
8'h63,
8'h73,
8'h3E,
8'h00,
8'h00,
8'h00,
8'h00,// 5
8'h00,
8'h00,
8'h1C,
8'h30,
8'h60,
8'h60,
8'h7E,
8'h63,
8'h63,
8'h63,
8'h63,
8'h3E,
8'h00,
8'h00,
8'h00,
8'h00,// 6
8'h00,
8'h00,
8'h7F,
8'h63,
8'h03,
8'h06,
8'h06,
8'h0C,
8'h0C,
8'h18,
8'h18,
8'h18,
8'h00,
8'h00,
8'h00,
8'h00,// 7
8'h00,
8'h00,
8'h3E,
8'h63,
8'h63,
8'h63,
8'h3E,
8'h63,
8'h63,
8'h63,
8'h63,
8'h3E,
8'h00,
8'h00,
8'h00,
8'h00,// 8
8'h00,
8'h00,
8'h3E,
8'h63,
8'h63,
8'h63,
8'h63,
8'h3F,
8'h03,
8'h03,
8'h06,
8'h3C,
8'h00,
8'h00,
8'h00,
8'h00,// 9
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h18,
8'h18,
8'h00,
8'h00,
8'h00,
8'h18,
8'h18,
8'h00,
8'h00,
8'h00,
8'h00,// :
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h18,
8'h18,
8'h00,
8'h00,
8'h00,
8'h18,
8'h18,
8'h18,
8'h30,
8'h00,
8'h00,// ;
8'h00,
8'h00,
8'h00,
8'h06,
8'h0C,
8'h18,
8'h30,
8'h60,
8'h30,
8'h18,
8'h0C,
8'h06,
8'h00,
8'h00,
8'h00,
8'h00,// <
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h7E,
8'h00,
8'h00,
8'h7E,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,// =
8'h00,
8'h00,
8'h00,
8'h60,
8'h30,
8'h18,
8'h0C,
8'h06,
8'h0C,
8'h18,
8'h30,
8'h60,
8'h00,
8'h00,
8'h00,
8'h00,// >
8'h00,
8'h00,
8'h3E,
8'h63,
8'h63,
8'h06,
8'h0C,
8'h0C,
8'h0C,
8'h00,
8'h0C,
8'h0C,
8'h00,
8'h00,
8'h00,
8'h00,// ?
8'h00,
8'h00,
8'h3E,
8'h63,
8'h63,
8'h6F,
8'h6B,
8'h6B,
8'h6E,
8'h60,
8'h60,
8'h3E,
8'h00,
8'h00,
8'h00,
8'h00,// @ 8'h40
8'h00,
8'h00,
8'h08,
8'h1C,
8'h36,
8'h63,
8'h63,
8'h63,
8'h7F,
8'h63,
8'h63,
8'h63,
8'h00,
8'h00,
8'h00,
8'h00,// A
8'h00,
8'h00,
8'h7E,
8'h33,
8'h33,
8'h33,
8'h3E,
8'h33,
8'h33,
8'h33,
8'h33,
8'h7E,
8'h00,
8'h00,
8'h00,
8'h00,// B
8'h00,
8'h00,
8'h1E,
8'h33,
8'h61,
8'h60,
8'h60,
8'h60,
8'h60,
8'h61,
8'h33,
8'h1E,
8'h00,
8'h00,
8'h00,
8'h00,// C
8'h00,
8'h00,
8'h7C,
8'h36,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h36,
8'h7C,
8'h00,
8'h00,
8'h00,
8'h00,// D
8'h00,
8'h00,
8'h7F,
8'h33,
8'h31,
8'h34,
8'h3C,
8'h34,
8'h30,
8'h31,
8'h33,
8'h7F,
8'h00,
8'h00,
8'h00,
8'h00,// E
8'h00,
8'h00,
8'h7F,
8'h33,
8'h31,
8'h34,
8'h3C,
8'h34,
8'h30,
8'h30,
8'h30,
8'h78,
8'h00,
8'h00,
8'h00,
8'h00,// F
8'h00,
8'h00,
8'h1E,
8'h33,
8'h61,
8'h60,
8'h60,
8'h6F,
8'h63,
8'h63,
8'h37,
8'h1D,
8'h00,
8'h00,
8'h00,
8'h00,// G
8'h00,
8'h00,
8'h63,
8'h63,
8'h63,
8'h63,
8'h7F,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h00,
8'h00,
8'h00,
8'h00,// H
8'h00,
8'h00,
8'h3C,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h3C,
8'h00,
8'h00,
8'h00,
8'h00,// I
8'h00,
8'h00,
8'h0F,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h66,
8'h66,
8'h3C,
8'h00,
8'h00,
8'h00,
8'h00,// J
8'h00,
8'h00,
8'h73,
8'h33,
8'h36,
8'h36,
8'h3C,
8'h36,
8'h36,
8'h33,
8'h33,
8'h73,
8'h00,
8'h00,
8'h00,
8'h00,// K
8'h00,
8'h00,
8'h78,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h31,
8'h33,
8'h7F,
8'h00,
8'h00,
8'h00,
8'h00,// L
8'h00,
8'h00,
8'h63,
8'h77,
8'h7F,
8'h6B,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h00,
8'h00,
8'h00,
8'h00,// M
8'h00,
8'h00,
8'h63,
8'h63,
8'h73,
8'h7B,
8'h7F,
8'h6F,
8'h67,
8'h63,
8'h63,
8'h63,
8'h00,
8'h00,
8'h00,
8'h00,// N
8'h00,
8'h00,
8'h1C,
8'h36,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h36,
8'h1C,
8'h00,
8'h00,
8'h00,
8'h00,// O
8'h00,
8'h00,
8'h7E,
8'h33,
8'h33,
8'h33,
8'h3E,
8'h30,
8'h30,
8'h30,
8'h30,
8'h78,
8'h00,
8'h00,
8'h00,
8'h00,// P   8'h50
8'h00,
8'h00,
8'h3E,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h6B,
8'h6F,
8'h3E,
8'h06,
8'h07,
8'h00,
8'h00,// Q
8'h00,
8'h00,
8'h7E,
8'h33,
8'h33,
8'h33,
8'h3E,
8'h36,
8'h36,
8'h33,
8'h33,
8'h73,
8'h00,
8'h00,
8'h00,
8'h00,// R
8'h00,
8'h00,
8'h3E,
8'h63,
8'h63,
8'h30,
8'h1C,
8'h06,
8'h03,
8'h63,
8'h63,
8'h3E,
8'h00,
8'h00,
8'h00,
8'h00,// S
8'h00,
8'h00,
8'hFF,
8'hDB,
8'h99,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h3C,
8'h00,
8'h00,
8'h00,
8'h00,// T
8'h00,
8'h00,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h3E,
8'h00,
8'h00,
8'h00,
8'h00,// U
8'h00,
8'h00,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h36,
8'h1C,
8'h08,
8'h00,
8'h00,
8'h00,
8'h00,// V
8'h00,
8'h00,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h6B,
8'h6B,
8'h7F,
8'h36,
8'h36,
8'h00,
8'h00,
8'h00,
8'h00,// W
8'h00,
8'h00,
8'hC3,
8'hC3,
8'h66,
8'h3C,
8'h18,
8'h18,
8'h3C,
8'h66,
8'hC3,
8'hC3,
8'h00,
8'h00,
8'h00,
8'h00,// X
8'h00,
8'h00,
8'hC3,
8'hC3,
8'hC3,
8'h66,
8'h3C,
8'h18,
8'h18,
8'h18,
8'h18,
8'h3C,
8'h00,
8'h00,
8'h00,
8'h00,// Y
8'h00,
8'h00,
8'h7F,
8'h63,
8'h43,
8'h06,
8'h0C,
8'h18,
8'h30,
8'h61,
8'h63,
8'h7F,
8'h00,
8'h00,
8'h00,
8'h00,// Z
8'h00,
8'h00,
8'h3C,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h30,
8'h3C,
8'h00,
8'h00,
8'h00,
8'h00,// [
8'h00,
8'h00,
8'h80,
8'hC0,
8'hE0,
8'h70,
8'h38,
8'h1C,
8'h0E,
8'h07,
8'h03,
8'h01,
8'h00,
8'h00,
8'h00,
8'h00,// \ (back slash)
8'h00,
8'h00,
8'h3C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h3C,
8'h00,
8'h00,
8'h00,
8'h00,// ]
8'h08,
8'h1C,
8'h36,
8'h63,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,// ^
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'hFF,
8'h00,
8'h00,
8'h00,// _
8'h18,
8'h18,
8'h0C,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,// `    8'h60
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h3C,
8'h46,
8'h06,
8'h3E,
8'h66,
8'h66,
8'h3B,
8'h00,
8'h00,
8'h00,
8'h00,// a
8'h00,
8'h00,
8'h70,
8'h30,
8'h30,
8'h3C,
8'h36,
8'h33,
8'h33,
8'h33,
8'h33,
8'h6E,
8'h00,
8'h00,
8'h00,
8'h00,// b
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h3E,
8'h63,
8'h60,
8'h60,
8'h60,
8'h63,
8'h3E,
8'h00,
8'h00,
8'h00,
8'h00,// c
8'h00,
8'h00,
8'h0E,
8'h06,
8'h06,
8'h1E,
8'h36,
8'h66,
8'h66,
8'h66,
8'h66,
8'h3B,
8'h00,
8'h00,
8'h00,
8'h00,// d
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h3E,
8'h63,
8'h63,
8'h7E,
8'h60,
8'h63,
8'h3E,
8'h00,
8'h00,
8'h00,
8'h00,// e
8'h00,
8'h00,
8'h1C,
8'h36,
8'h32,
8'h30,
8'h7C,
8'h30,
8'h30,
8'h30,
8'h30,
8'h78,
8'h00,
8'h00,
8'h00,
8'h00,// f
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h3B,
8'h66,
8'h66,
8'h66,
8'h66,
8'h3E,
8'h06,
8'h66,
8'h3C,
8'h00,
8'h00,// g
8'h00,
8'h00,
8'h70,
8'h30,
8'h30,
8'h36,
8'h3B,
8'h33,
8'h33,
8'h33,
8'h33,
8'h73,
8'h00,
8'h00,
8'h00,
8'h00,// h
8'h00,
8'h00,
8'h0C,
8'h0C,
8'h00,
8'h1C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h1E,
8'h00,
8'h00,
8'h00,
8'h00,// i
8'h00,
8'h00,
8'h06,
8'h06,
8'h00,
8'h0E,
8'h06,
8'h06,
8'h06,
8'h06,
8'h06,
8'h66,
8'h66,
8'h3C,
8'h00,
8'h00,// j
8'h00,
8'h00,
8'h70,
8'h30,
8'h30,
8'h33,
8'h33,
8'h36,
8'h3C,
8'h36,
8'h33,
8'h73,
8'h00,
8'h00,
8'h00,
8'h00,// k
8'h00,
8'h00,
8'h1C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h0C,
8'h1E,
8'h00,
8'h00,
8'h00,
8'h00,// l
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h6E,
8'h7F,
8'h6B,
8'h6B,
8'h6B,
8'h6B,
8'h6B,
8'h00,
8'h00,
8'h00,
8'h00,// m
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h6E,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h33,
8'h00,
8'h00,
8'h00,
8'h00,// n
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h3E,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h3E,
8'h00,
8'h00,
8'h00,
8'h00,// o
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h6E,
8'h33,
8'h33,
8'h33,
8'h33,
8'h3E,
8'h30,
8'h30,
8'h78,
8'h00,
8'h00,// p    8'h70
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h3B,
8'h66,
8'h66,
8'h66,
8'h66,
8'h3E,
8'h06,
8'h06,
8'h0F,
8'h00,
8'h00,// q
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h6E,
8'h3B,
8'h33,
8'h30,
8'h30,
8'h30,
8'h78,
8'h00,
8'h00,
8'h00,
8'h00,// r
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h3E,
8'h63,
8'h38,
8'h0E,
8'h03,
8'h63,
8'h3E,
8'h00,
8'h00,
8'h00,
8'h00,// s
8'h00,
8'h00,
8'h08,
8'h18,
8'h18,
8'h7E,
8'h18,
8'h18,
8'h18,
8'h18,
8'h1B,
8'h0E,
8'h00,
8'h00,
8'h00,
8'h00,// t
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h66,
8'h66,
8'h66,
8'h66,
8'h66,
8'h66,
8'h3B,
8'h00,
8'h00,
8'h00,
8'h00,// u
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h63,
8'h63,
8'h36,
8'h36,
8'h1C,
8'h1C,
8'h08,
8'h00,
8'h00,
8'h00,
8'h00,// v
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h63,
8'h63,
8'h63,
8'h6B,
8'h6B,
8'h7F,
8'h36,
8'h00,
8'h00,
8'h00,
8'h00,// w
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h63,
8'h36,
8'h1C,
8'h1C,
8'h1C,
8'h36,
8'h63,
8'h00,
8'h00,
8'h00,
8'h00,// x
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h63,
8'h63,
8'h63,
8'h63,
8'h63,
8'h3F,
8'h03,
8'h06,
8'h3C,
8'h00,
8'h00,// y
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h7F,
8'h66,
8'h0C,
8'h18,
8'h30,
8'h63,
8'h7F,
8'h00,
8'h00,
8'h00,
8'h00,// z
8'h00,
8'h00,
8'h0E,
8'h18,
8'h18,
8'h18,
8'h70,
8'h18,
8'h18,
8'h18,
8'h18,
8'h0E,
8'h00,
8'h00,
8'h00,
8'h00,// 
8'h00,
8'h00,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h00,
8'h18,
8'h18,
8'h18,
8'h18,
8'h18,
8'h00,
8'h00,
8'h00,// |
8'h00,
8'h00,
8'h70,
8'h18,
8'h18,
8'h18,
8'h0E,
8'h18,
8'h18,
8'h18,
8'h18,
8'h70,
8'h00,
8'h00,
8'h00,
8'h00,// }
8'h00,
8'h00,
8'h3B,
8'h6E,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,// ~
8'h00,
8'h70,
8'hD8,
8'hD8,
8'h70,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00,
8'h00 // DEL
};