parameter [0:7] char_rom_y [0:159] = {
8'b00000000,
8'b00000000,
8'b00011000,
8'b00111000,
8'b01111000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b01111110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01111100,
8'b11000110,
8'b00000110,
8'b00001100,
8'b00011000,
8'b00110000,
8'b01100000,
8'b11000000,
8'b11000110,
8'b11111110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01111100,
8'b11000110,
8'b00000110,
8'b00000110,
8'b00111100,
8'b00000110,
8'b00000110,
8'b00000110,
8'b11000110,
8'b01111100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00001100,
8'b00011100,
8'b00111100,
8'b01101100,
8'b11001100,
8'b11111110,
8'b00001100,
8'b00001100,
8'b00001100,
8'b00011110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b11111110,
8'b11000000,
8'b11000000,
8'b11000000,
8'b11111100,
8'b00000110,
8'b00000110,
8'b00000110,
8'b11000110,
8'b01111100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111000,
8'b01100000,
8'b11000000,
8'b11000000,
8'b11111100,
8'b11000110,
8'b11000110,
8'b11000110,
8'b11000110,
8'b01111100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b11111110,
8'b11000110,
8'b00000110,
8'b00000110,
8'b00001100,
8'b00011000,
8'b00110000,
8'b00110000,
8'b00110000,
8'b00110000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01111100,
8'b11000110,
8'b11000110,
8'b11000110,
8'b01111100,
8'b11000110,
8'b11000110,
8'b11000110,
8'b11000110,
8'b01111100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01111100,
8'b11000110,
8'b11000110,
8'b11000110,
8'b01111110,
8'b00000110,
8'b00000110,
8'b00000110,
8'b00001100,
8'b01111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01111100,
8'b11000110,
8'b11000110,
8'b11001110,
8'b11011110,
8'b11110110,
8'b11100110,
8'b11000110,
8'b11000110,
8'b01111100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000
};
