parameter [0:7] char_rom_x [0:303] = {
8'b00000000,
8'b00000000,
8'b00010000,
8'b00111000,
8'b01101100,
8'b11000110,
8'b11000110,
8'b11111110,
8'b11000110,
8'b11000110,
8'b11000110,
8'b11000110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b11111100,
8'b01100110,
8'b01100110,
8'b01100110,
8'b01111100,
8'b01100110,
8'b01100110,
8'b01100110,
8'b01100110,
8'b11111100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111100,
8'b01100110,
8'b11000010,
8'b11000000,
8'b11000000,
8'b11000000,
8'b11000000,
8'b11000010,
8'b01100110,
8'b00111100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b11111000,
8'b01101100,
8'b01100110,
8'b01100110,
8'b01100110,
8'b01100110,
8'b01100110,
8'b01100110,
8'b01101100,
8'b11111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b11111110,
8'b01100110,
8'b01100010,
8'b01101000,
8'b01111000,
8'b01101000,
8'b01100000,
8'b01100010,
8'b01100110,
8'b11111110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b11111110,
8'b01100110,
8'b01100010,
8'b01101000,
8'b01111000,
8'b01101000,
8'b01100000,
8'b01100000,
8'b01100000,
8'b11110000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111100,
8'b01100110,
8'b11000010,
8'b11000000,
8'b11000000,
8'b11011110,
8'b11000110,
8'b11000110,
8'b01100110,
8'b00111010,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b11000110,
8'b11000110,
8'b11000110,
8'b11000110,
8'b11111110,
8'b11000110,
8'b11000110,
8'b11000110,
8'b11000110,
8'b11000110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00011110,
8'b00001100,
8'b00001100,
8'b00001100,
8'b00001100,
8'b00001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b01111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b11100110,
8'b01100110,
8'b01100110,
8'b01101100,
8'b01111000,
8'b01111000,
8'b01101100,
8'b01100110,
8'b01100110,
8'b11100110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b11110000,
8'b01100000,
8'b01100000,
8'b01100000,
8'b01100000,
8'b01100000,
8'b01100000,
8'b01100010,
8'b01100110,
8'b11111110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b11000011,
8'b11100111,
8'b11111111,
8'b11111111,
8'b11011011,
8'b11000011,
8'b11000011,
8'b11000011,
8'b11000011,
8'b11000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b11000110,
8'b11100110,
8'b11110110,
8'b11111110,
8'b11011110,
8'b11001110,
8'b11000110,
8'b11000110,
8'b11000110,
8'b11000110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01111100,
8'b11000110,
8'b11000110,
8'b11000110,
8'b11000110,
8'b11000110,
8'b11000110,
8'b11000110,
8'b11000110,
8'b01111100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b11111100,
8'b01100110,
8'b01100110,
8'b01100110,
8'b01111100,
8'b01100000,
8'b01100000,
8'b01100000,
8'b01100000,
8'b11110000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01111100,
8'b11000110,
8'b11000110,
8'b11000110,
8'b11000110,
8'b11000110,
8'b11000110,
8'b11010110,
8'b11011110,
8'b01111100,
8'b00001100,
8'b00001110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b11111100,
8'b01100110,
8'b01100110,
8'b01100110,
8'b01111100,
8'b01101100,
8'b01100110,
8'b01100110,
8'b01100110,
8'b11100110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01111100,
8'b11000110,
8'b11000110,
8'b01100000,
8'b00111000,
8'b00001100,
8'b00000110,
8'b11000110,
8'b11000110,
8'b01111100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b11111111,
8'b11011011,
8'b10011001,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00011000,
8'b00111100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000
};
